package i2c_pkg;
    import ncsu_pkg::*;
    /* `include "ncsu_macros.svh" */
    `include "../../ncsu_pkg/ncsu_macros.svh"

    `include "src/i2c_typedefs.svh"
    `include "src/i2c_configuration.svh"
    `include "src/i2c_transaction_base.svh"
    `include "src/i2c_driver.svh"
    `include "src/i2c_monitor.svh"
    /* `include "src/i2c_coverage.svh" */
    `include "src/i2c_agent.svh"
    /* `include "src/i2c_if.sv" */

endpackage
