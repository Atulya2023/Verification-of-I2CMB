typedef enum bit [1:0] {CSR, DPR, CMDR, FSM} wb_reg;
typedef enum bit {WRITE, READ} wb_op_t;
