typedef enum bit {WRITE_OP, READ_OP} i2c_op_t;
