class i2cmb_test extends generator;
    `ncsu_register_object(i2cmb_test)
endclass
